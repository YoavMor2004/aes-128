module sub_bytes (
    input  logic [127:0] in_bus,   // 128-bit input bus
    output logic [127:0] out_bus   // 128-bit output bus
);

    // Module logic goes here

endmodule
