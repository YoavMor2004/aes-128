module sbox (
    input  logic [7:0] in_bus,   // 8-bit input bus
    output logic [7:0] out_bus   // 8-bit output bus
);

    // Module logic goes here

endmodule
